module top;
   import uvm_pkg::*;
`include "uvm_macros.svh"

   import example_pkg::*;

   initial run_test("communication_test");
endmodule : top

     