   typedef struct {
      byte unsigned        A;
      byte unsigned        B;
      operation_t op;
   } command_s;