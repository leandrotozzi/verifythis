package dice_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   
   `include "dice_roller.svh"       
   `include "coverage.svh"
   `include "histogram.svh"
   `include "average.svh"
   `include "dice_test.svh"
   
endpackage : dice_pkg
   
   