module top;
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   import dice_pkg::*;
   initial run_test("dice_test");
endmodule : top

