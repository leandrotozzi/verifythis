   // Constructor para uvm_object. Ultra Sencillo
   function new (string name = "");
      super.new(name);
   endfunction : new